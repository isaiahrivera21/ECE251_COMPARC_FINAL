////////////////////////////////////////////////////////////////////////////////
//      
//      Module: module_name 
//      Hdl: Verilog
//
//      Module Description: 
//
//      Author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef EXAMPLE
`define EXAMPLE

module example();

   //
   // ---------------- PARAMETER DECLARATIONS ----------------
   //

   //
   // ---------------- PORT DEFINITIONS ----------------
   //


   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //


endmodule

`endif // EXAMPLE

